module mult

endmodule