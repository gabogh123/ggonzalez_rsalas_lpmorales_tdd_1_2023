module current_state_new_tile_check();



endmodule
