module new_tile_check_tb();



endmodule
