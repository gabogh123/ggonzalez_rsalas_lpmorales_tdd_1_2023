/*

Extend

*/
module extend
    #  (parameter N = 24)
	   (A, S, Y);

    input  logic [N-1:0] A;
    input  logic         S;
	output logic  [31:0] Y;



endmodule