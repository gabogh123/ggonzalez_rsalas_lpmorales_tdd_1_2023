module next_state_new_tile_check();




endmodule
