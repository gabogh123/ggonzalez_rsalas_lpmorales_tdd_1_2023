/*
Test Bench para MUX 32:1 parametrizable para N bits
*/
module mux32NtoN_tb;

	parameter integer N = 32;

	logic [N-1:0] I00;
    logic [N-1:0] I01;
    logic [N-1:0] I02;
    logic [N-1:0] I03;
    logic [N-1:0] I04;
    logic [N-1:0] I05;
    logic [N-1:0] I06;
    logic [N-1:0] I07;
    logic [N-1:0] I08;
    logic [N-1:0] I09;
    logic [N-1:0] I10; 
    logic [N-1:0] I11;
    logic [N-1:0] I12;
    logic [N-1:0] I13;
    logic [N-1:0] I14;
    logic [N-1:0] I15;
    logic [N-1:0] I16;
    logic [N-1:0] I17;
    logic [N-1:0] I18;
    logic [N-1:0] I19;
    logic [N-1:0] I20;
    logic [N-1:0] I21;
    logic [N-1:0] I22;
    logic [N-1:0] I23;
    logic [N-1:0] I24;
    logic [N-1:0] I25;
    logic [N-1:0] I26;
    logic [N-1:0] I27;
    logic [N-1:0] I28;
    logic [N-1:0] I29;
    logic [N-1:0] I30;
    logic [N-1:0] I31;

	logic    [4:0]  S;
	logic      enable;
	logic  [N-1:0]  O;	

	mux_32NtoN # (.N(N)) uut (.I00(I00),
							  .I01(I01),
							  .I02(I02),
							  .I03(I03),
							  .I04(I04),
							  .I05(I05),
							  .I06(I06),
							  .I07(I07),
							  .I08(I08),
							  .I09(I09),
							  .I10(I10),
							  .I11(I11),
							  .I12(I12),
							  .I13(I13),
							  .I14(I14),
							  .I15(I15),
							  .I16(I16),
							  .I17(I17),
							  .I18(I18),
							  .I19(I19),
							  .I20(I20),
							  .I21(I21),
							  .I22(I22),
							  .I23(I23),
							  .I24(I24),
							  .I25(I25),
							  .I26(I26),
							  .I27(I27),
							  .I28(I28),
							  .I29(I29),
							  .I30(I30),
							  .I31(I31),
							  .S(S),
							  .enable(enable),
							  .O(O));

	initial begin
		$display("mux32NtoN Test Bench:\n");

		I00 <= 32'b0;
		I01 <= 32'b0;
		I02 <= 32'b0;
		I03 <= 32'b0;
		I04 <= 32'b0;
		I05 <= 32'b0;
		I06 <= 32'b0;
		I07 <= 32'b0;
		I08 <= 32'b0;
		I09 <= 32'b0;
		I10 <= 32'b0;
		I11 <= 32'b0;
		I12 <= 32'b0;
		I13 <= 32'b0;
		I14 <= 32'b0;
		I15 <= 32'b0;
		I16 <= 32'b0;
		I17 <= 32'b0;
		I18 <= 32'b0;
		I19 <= 32'b0;
		I20 <= 32'b0;
		I21 <= 32'b0;
		I22 <= 32'b0;
		I23 <= 32'b0;
		I24 <= 32'b0;
		I25 <= 32'b0;
		I26 <= 32'b0;
		I27 <= 32'b0;
		I28 <= 32'b0;
		I29 <= 32'b0;
		I30 <= 32'b0;
		I31 <= 32'b0;
		
		S <= 5'b00000;
		enable <= 0;

		$monitor("S=%b enable=%b\n", S, enable,
				 "I00=%b I01=%b I02=%b I03=%b\n", I00, I01, I02, I03,
				 "I04=%b I05=%b I06=%b I07=%b\n", I04, I05, I06, I07,
				 "I08=%b I09=%b I10=%b I11=%b\n", I08, I09, I10, I11,
				 "I12=%b I13=%b I14=%b I15=%b\n", I12, I13, I14, I15,
				 "I16=%b I17=%b I18=%b I19=%b\n", I16, I17, I18, I19,
				 "I20=%b I21=%b I22=%b I23=%b\n", I20, I21, I22, I23,
				 "I24=%b I25=%b I26=%b I27=%b\n", I24, I25, I26, I27,
				 "I28=%b I29=%b I30=%b I31=%b\n", I28, I29, I30, I31,
				 "O=%b\n", O);
	end

	initial	begin
	
		#100

        enable = 1;

        #100

		I00 <= 32'b11100101100111110001000000100000;
		I01 <= 32'b10101010000000000000000000000100;
		I02 <= 32'b11100011101000000000000000000000;
		I03 <= 32'b11100001101000000010000010100010;
		I04 <= 32'b11101000100101011101001001110101;
		I05 <= 32'b01010000000010101001110101001001;
		I06 <= 32'b00010010001000100010010110101000;
		I07 <= 32'b11111010110110110110111011011011;
		I08 <= 32'b00101000101001000100111010101111;
		I09 <= 32'b01010010001001001001000100101010;
		I10 <= 32'b11101010101011111101000000100000;
		I11 <= 32'b10101010001111110110111100000100;
		I12 <= 32'b11100011101000101010010111010100;
		I13 <= 32'b11100001101000001011010110010010;
		I14 <= 32'b01001000101010101011101001110101;
		I15 <= 32'b01010010101101101011110101001001;
		I16 <= 32'b00010010001010011010010101111010;
		I17 <= 32'b11111010000000110101110110011011;
		I18 <= 32'b00101000101001110101101010000011;
		I19 <= 32'b01010101011110001001000100101010;
		I20 <= 32'b11101010101000010010101010000000;
		I21 <= 32'b10101010000000010011011111111110;
		I22 <= 32'b11100000101010101111101010010100;
		I23 <= 32'b00101001011100101011010110010010;
		I24 <= 32'b01010101001111111011101001110101;
		I25 <= 32'b01010010111010100000101011001001;
		I26 <= 32'b00010010001000000101101110101000;
		I27 <= 32'b10100101010101111010010110011011;
		I28 <= 32'b00101000000010101011101010000011;
		I29 <= 32'b11111010101000001001000100101010;
		I30 <= 32'b11101010000101010111111111110000;
		I31 <= 32'b010111111101010001000101011001001;

		#100

		S <= 5'b00000;

        #100

        // assert

        #100

        S <= 5'b00010;

        #100

        // assert

        #100

        S <= 5'b01010;

        #100

        // assert

        #100

        enable = 0;

        #100

        S <= 5'b11110;

        #100

        // assert

        #100

        S <= 5'b10110;

        #100

        // assert

		#100;

        // Done

    end

endmodule
