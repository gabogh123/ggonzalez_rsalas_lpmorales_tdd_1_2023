module alu_p_tb;

    parameter integer N = 32;

    logic [N-1:0]     A;
	logic [N-1:0]     B;
	logic   [3:0]  func;
	logic [N-1:0]     Y;
	logic   [3:0] flags;

    alu # (.N(N)) uut (.A(A),
                       .B(B),
                       .func(func),
                       .Y(Y),
                       .flags(flags));

    initial begin
		$display("alu Test Bench:\n");

		A = 0;
        B = 0;
        func = 0;

		$monitor("func: %b\nA = %b *func* B = %b\nY = %b\nflags: %b\n",
                 func, A, B, Y, flags);

	end

    initial	begin

		#200

        $display("0. 0000 = sum:\n");
        A <= 32'b11100101100111110001000000100000;
		B <= 32'b00000000000000000000000000000100;
        func = 4'b0000;

        #100
        	
		assert((Y === 32'b11100101100111110001000000100100) & (flags === 4'b0000))
        else $error("Failed");
	
		#100

        $display("1. 0001 = sub:\n");
        A <= 32'b11100101100111110001000000100101;
		B <= 32'b00000000000000000000000000000100;
        func = 4'b0001;

        #100
        	
		assert((Y === 32'b11100101100111110001000000100001) & (flags === 4'b0000))
        else $error("Failed");

        #100

        $display("2. 0010 = mult:\n");
        A <= 32'b00000000000001010100101001001001;
		B <= 32'b00000000000000000010001001011101;
        func = 4'b0010;

        #100
        	
		assert((Y === 32'b10110101110010011010111010000101) & (flags === 4'b0000))
        else $error("Failed");

        #100
        /*
        $display("3. 0011 = div:\n");
        A <= 32'b01000010001010110101101111101010;
		B <= 32'b00001001000010000101000101010101;
        func = 4'b0011;
        
        #100
        	
		assert((Y === 32'b00000010111100010010001010010111) & (flags === 4'b0000))
        else $error("Failed");
        */
        #100
        /*
        $display("4. 0100 = mod:\n");
        A <= 32'b10111001000111001000100001110011;
		B <= 32'b00100000101011110101100100010100;
        func = 4'b0100;
        
        #100
        	
		assert((Y === 32'b00010101101011111100101100001111) & (flags === 4'b0000))
        else $error("Failed");
        */
        #100

        $display("5. 0101 = and:\n");
        A <= 32'b11101011101000101101110001001010;
		B <= 32'b01001010101011101010101010010101;
        func = 4'b0101;

        #100
        	
		assert((Y === 32'b01001010101000101000100000000000) & (flags === 4'b0000))
        else $error("Failed");

        #100

        $display("6. 0110 = or:\n");
        A <= 32'b01101011101000101101110001001010;
		B <= 32'b00100101010100100101001001000101;
        func = 4'b0110;

        #100
        	
		assert((Y === 32'b01101111111100101101111001001111) & (flags === 4'b0000))
        else $error("Failed");

        #100

        $display("7. 0111 = xor:\n");
        A <= 32'b00101010011011001010101001011000;
		B <= 32'b10010101001010101101001011111101;
                
        func = 4'b0111;

        #100
        	
		assert((Y === 32'b10111111010001100111100010100101) & (flags === 4'b0000))
        else $error("Failed");

        #100
        /*
        $display("8. 1000 = shift L:\n");
        A <= 32'b10100101001010011101010101001010;
		B <= 32'b00000000000000000000000000000001;
        func = 4'b1000;

        #100
        	
		assert((Y === 32'b0) & (flags === 4'b0000))
        else $error("Failed");
        */
        #100
        /*
        $display("9. 1001 = shift R:\n");
        A <= 32'b01001000001010100101010110101010;
		B <= 32'b00000000000000000000000000000011;
        func = 4'b1001;

        #100
        	
		assert((Y === 32'b0) & (flags === 4'b0000))
        else $error("Failed");
        */
		#100;

        // Semidone

    end

endmodule