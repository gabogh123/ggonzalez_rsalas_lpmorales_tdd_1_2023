module resta


endmodule