/*

ALU

*/
module alu(A, B, func, Y, flags);

    input  [31:0]     A;
    input  [31:0]     B;
    input   [3:0]  func;
    output [31:0]     Y;
    output  [4:0] flags;


endmodule