module div

endmodule