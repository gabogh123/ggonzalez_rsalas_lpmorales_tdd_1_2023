module histogram_equalizer(A, B);

	input  logic A;
	output logic B;

endmodule