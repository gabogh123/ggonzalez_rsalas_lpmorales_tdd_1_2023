module resta(a,b,y,c);




endmodule