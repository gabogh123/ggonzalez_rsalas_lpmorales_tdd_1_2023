
module histogram_equalizer_tb;

	

endmodule
